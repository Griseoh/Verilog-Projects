$date
	Sun Sep 24 05:14:32 2023
$end
$version
	Icarus Verilog
$end
$timescale
	1ns
$end
$scope module Comparator_2bit_tb $end
$var wire 6 ! Y [5:0] $end
$var reg 2 " A [1:0] $end
$var reg 2 # B [1:0] $end
$scope module uut $end
$var wire 2 $ A [1:0] $end
$var wire 2 % B [1:0] $end
$var reg 6 & Y [5:0] $end
$upscope $end
$upscope $end
$enddefinitions $end
$comment Show the parameter values. $end
$dumpall
$end
#0
$dumpvars
bx &
bx %
bx $
bx #
bx "
bx !
$end
#5
b100011 !
b100011 &
b0 #
b0 %
b0 "
b0 $
#10
b10101 !
b10101 &
b1 #
b1 %
#15
b10 #
b10 %
#20
b11 #
b11 %
#25
b11010 !
b11010 &
b0 #
b0 %
b1 "
b1 $
#30
b100011 !
b100011 &
b1 #
b1 %
#35
b10101 !
b10101 &
b10 #
b10 %
#40
b11 #
b11 %
#45
b11010 !
b11010 &
b0 #
b0 %
b10 "
b10 $
#50
b1 #
b1 %
#55
b100011 !
b100011 &
b10 #
b10 %
#60
b10101 !
b10101 &
b11 #
b11 %
#65
b11010 !
b11010 &
b0 #
b0 %
b11 "
b11 $
#70
b1 #
b1 %
#75
b10 #
b10 %
#80
b100011 !
b100011 &
b11 #
b11 %
#90
