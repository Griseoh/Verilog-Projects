module simpleand (f, a, b);
    input a,b;
    output f;
    assign f = a&b;
endmodule